`default_nettype none

// module mul4
//    (  input wire [3:0]  x1,
//       input wire [3:0]  x2,
//       output wire [7:0] y);

//    assign y = (x1 == 4'b0) ? {8'b0} :
//               (x2 == 4'b0) ? {8'b0} :
//               (x1 == 4'b1) ? {4'b0,x2} :
//               (x2 == 4'b1) ? {4'b0,x1} :
//               (x1 == 4'b10) ? {3'b0,x2,1'b0} :
//               (x2 == 4'b10) ? {3'b0,x1,1'b0} :
//               (x1 == 4'b100) ? {2'b0,x2,2'b0} :
//               (x2 == 4'b100) ? {2'b0,x1,2'b0} :
//               (x1 == 4'b1000) ? {1'b0,x2,3'b0} :
//               (x2 == 4'b1000) ? {1'b0,x1,3'b0} :
//               (x1 == 4'b11 && x2 == 4'b11) ? {8'b1001} :
//               (x1 == 4'b11 && x2 == 4'b101) ? {8'b1111} :
//               (x1 == 4'b11 && x2 == 4'b110) ? {8'b10010} :
//               (x1 == 4'b11 && x2 == 4'b111) ? {8'b10101} :
//               (x1 == 4'b11 && x2 == 4'b1001) ? {8'b11011} :
//               (x1 == 4'b11 && x2 == 4'b1010) ? {8'b11110} :
//               (x1 == 4'b11 && x2 == 4'b1011) ? {8'b100001} :
//               (x1 == 4'b11 && x2 == 4'b1100) ? {8'b100100} :
//               (x1 == 4'b11 && x2 == 4'b1101) ? {8'b100111} :
//               (x1 == 4'b11 && x2 == 4'b1110) ? {8'b101010} :
//               (x1 == 4'b11 && x2 == 4'b1111) ? {8'b101101} :
//               (x1 == 4'b101 && x2 == 4'b11) ? {8'b1111} :
//               (x1 == 4'b101 && x2 == 4'b101) ? {8'b11001} :
//               (x1 == 4'b101 && x2 == 4'b110) ? {8'b11110} :
//               (x1 == 4'b101 && x2 == 4'b111) ? {8'b100011} :
//               (x1 == 4'b101 && x2 == 4'b1001) ? {8'b101101} :
//               (x1 == 4'b101 && x2 == 4'b1010) ? {8'b110010} :
//               (x1 == 4'b101 && x2 == 4'b1011) ? {8'b110111} :
//               (x1 == 4'b101 && x2 == 4'b1100) ? {8'b111100} :
//               (x1 == 4'b101 && x2 == 4'b1101) ? {8'b1000001} :
//               (x1 == 4'b101 && x2 == 4'b1110) ? {8'b1000110} :
//               (x1 == 4'b101 && x2 == 4'b1111) ? {8'b1001011} :
//               (x1 == 4'b110 && x2 == 4'b11) ? {8'b10010} :
//               (x1 == 4'b110 && x2 == 4'b101) ? {8'b11110} :
//               (x1 == 4'b110 && x2 == 4'b110) ? {8'b100100} :
//               (x1 == 4'b110 && x2 == 4'b111) ? {8'b101010} :
//               (x1 == 4'b110 && x2 == 4'b1001) ? {8'b110110} :
//               (x1 == 4'b110 && x2 == 4'b1010) ? {8'b111100} :
//               (x1 == 4'b110 && x2 == 4'b1011) ? {8'b1000010} :
//               (x1 == 4'b110 && x2 == 4'b1100) ? {8'b1001000} :
//               (x1 == 4'b110 && x2 == 4'b1101) ? {8'b1001110} :
//               (x1 == 4'b110 && x2 == 4'b1110) ? {8'b1010100} :
//               (x1 == 4'b110 && x2 == 4'b1111) ? {8'b1011010} :
//               (x1 == 4'b111 && x2 == 4'b11) ? {8'b10101} :
//               (x1 == 4'b111 && x2 == 4'b101) ? {8'b100011} :
//               (x1 == 4'b111 && x2 == 4'b110) ? {8'b101010} :
//               (x1 == 4'b111 && x2 == 4'b111) ? {8'b110001} :
//               (x1 == 4'b111 && x2 == 4'b1001) ? {8'b111111} :
//               (x1 == 4'b111 && x2 == 4'b1010) ? {8'b1000110} :
//               (x1 == 4'b111 && x2 == 4'b1011) ? {8'b1001101} :
//               (x1 == 4'b111 && x2 == 4'b1100) ? {8'b1010100} :
//               (x1 == 4'b111 && x2 == 4'b1101) ? {8'b1011011} :
//               (x1 == 4'b111 && x2 == 4'b1110) ? {8'b1100010} :
//               (x1 == 4'b111 && x2 == 4'b1111) ? {8'b1101001} :
//               (x1 == 4'b1001 && x2 == 4'b11) ? {8'b11011} :
//               (x1 == 4'b1001 && x2 == 4'b101) ? {8'b101101} :
//               (x1 == 4'b1001 && x2 == 4'b110) ? {8'b110110} :
//               (x1 == 4'b1001 && x2 == 4'b111) ? {8'b111111} :
//               (x1 == 4'b1001 && x2 == 4'b1001) ? {8'b1010001} :
//               (x1 == 4'b1001 && x2 == 4'b1010) ? {8'b1011010} :
//               (x1 == 4'b1001 && x2 == 4'b1011) ? {8'b1100011} :
//               (x1 == 4'b1001 && x2 == 4'b1100) ? {8'b1101100} :
//               (x1 == 4'b1001 && x2 == 4'b1101) ? {8'b1110101} :
//               (x1 == 4'b1001 && x2 == 4'b1110) ? {8'b1111110} :
//               (x1 == 4'b1001 && x2 == 4'b1111) ? {8'b10000111} :
//               (x1 == 4'b1010 && x2 == 4'b11) ? {8'b11110} :
//               (x1 == 4'b1010 && x2 == 4'b101) ? {8'b110010} :
//               (x1 == 4'b1010 && x2 == 4'b110) ? {8'b111100} :
//               (x1 == 4'b1010 && x2 == 4'b111) ? {8'b1000110} :
//               (x1 == 4'b1010 && x2 == 4'b1001) ? {8'b1011010} :
//               (x1 == 4'b1010 && x2 == 4'b1010) ? {8'b1100100} :
//               (x1 == 4'b1010 && x2 == 4'b1011) ? {8'b1101110} :
//               (x1 == 4'b1010 && x2 == 4'b1100) ? {8'b1111000} :
//               (x1 == 4'b1010 && x2 == 4'b1101) ? {8'b10000010} :
//               (x1 == 4'b1010 && x2 == 4'b1110) ? {8'b10001100} :
//               (x1 == 4'b1010 && x2 == 4'b1111) ? {8'b10010110} :
//               (x1 == 4'b1011 && x2 == 4'b11) ? {8'b100001} :
//               (x1 == 4'b1011 && x2 == 4'b101) ? {8'b110111} :
//               (x1 == 4'b1011 && x2 == 4'b110) ? {8'b1000010} :
//               (x1 == 4'b1011 && x2 == 4'b111) ? {8'b1001101} :
//               (x1 == 4'b1011 && x2 == 4'b1001) ? {8'b1100011} :
//               (x1 == 4'b1011 && x2 == 4'b1010) ? {8'b1101110} :
//               (x1 == 4'b1011 && x2 == 4'b1011) ? {8'b1111001} :
//               (x1 == 4'b1011 && x2 == 4'b1100) ? {8'b10000100} :
//               (x1 == 4'b1011 && x2 == 4'b1101) ? {8'b10001111} :
//               (x1 == 4'b1011 && x2 == 4'b1110) ? {8'b10011010} :
//               (x1 == 4'b1011 && x2 == 4'b1111) ? {8'b10100101} :
//               (x1 == 4'b1100 && x2 == 4'b11) ? {8'b100100} :
//               (x1 == 4'b1100 && x2 == 4'b101) ? {8'b111100} :
//               (x1 == 4'b1100 && x2 == 4'b110) ? {8'b1001000} :
//               (x1 == 4'b1100 && x2 == 4'b111) ? {8'b1010100} :
//               (x1 == 4'b1100 && x2 == 4'b1001) ? {8'b1101100} :
//               (x1 == 4'b1100 && x2 == 4'b1010) ? {8'b1111000} :
//               (x1 == 4'b1100 && x2 == 4'b1011) ? {8'b10000100} :
//               (x1 == 4'b1100 && x2 == 4'b1100) ? {8'b10010000} :
//               (x1 == 4'b1100 && x2 == 4'b1101) ? {8'b10011100} :
//               (x1 == 4'b1100 && x2 == 4'b1110) ? {8'b10101000} :
//               (x1 == 4'b1100 && x2 == 4'b1111) ? {8'b10110100} :
//               (x1 == 4'b1101 && x2 == 4'b11) ? {8'b100111} :
//               (x1 == 4'b1101 && x2 == 4'b101) ? {8'b1000001} :
//               (x1 == 4'b1101 && x2 == 4'b110) ? {8'b1001110} :
//               (x1 == 4'b1101 && x2 == 4'b111) ? {8'b1011011} :
//               (x1 == 4'b1101 && x2 == 4'b1001) ? {8'b1110101} :
//               (x1 == 4'b1101 && x2 == 4'b1010) ? {8'b10000010} :
//               (x1 == 4'b1101 && x2 == 4'b1011) ? {8'b10001111} :
//               (x1 == 4'b1101 && x2 == 4'b1100) ? {8'b10011100} :
//               (x1 == 4'b1101 && x2 == 4'b1101) ? {8'b10101001} :
//               (x1 == 4'b1101 && x2 == 4'b1110) ? {8'b10110110} :
//               (x1 == 4'b1101 && x2 == 4'b1111) ? {8'b11000011} :
//               (x1 == 4'b1110 && x2 == 4'b11) ? {8'b101010} :
//               (x1 == 4'b1110 && x2 == 4'b101) ? {8'b1000110} :
//               (x1 == 4'b1110 && x2 == 4'b110) ? {8'b1010100} :
//               (x1 == 4'b1110 && x2 == 4'b111) ? {8'b1100010} :
//               (x1 == 4'b1110 && x2 == 4'b1001) ? {8'b1111110} :
//               (x1 == 4'b1110 && x2 == 4'b1010) ? {8'b10001100} :
//               (x1 == 4'b1110 && x2 == 4'b1011) ? {8'b10011010} :
//               (x1 == 4'b1110 && x2 == 4'b1100) ? {8'b10101000} :
//               (x1 == 4'b1110 && x2 == 4'b1101) ? {8'b10110110} :
//               (x1 == 4'b1110 && x2 == 4'b1110) ? {8'b11000100} :
//               (x1 == 4'b1110 && x2 == 4'b1111) ? {8'b11010010} :
//               (x1 == 4'b1111 && x2 == 4'b11) ? {8'b101101} :
//               (x1 == 4'b1111 && x2 == 4'b101) ? {8'b1001011} :
//               (x1 == 4'b1111 && x2 == 4'b110) ? {8'b1011010} :
//               (x1 == 4'b1111 && x2 == 4'b111) ? {8'b1101001} :
//               (x1 == 4'b1111 && x2 == 4'b1001) ? {8'b10000111} :
//               (x1 == 4'b1111 && x2 == 4'b1010) ? {8'b10010110} :
//               (x1 == 4'b1111 && x2 == 4'b1011) ? {8'b10100101} :
//               (x1 == 4'b1111 && x2 == 4'b1100) ? {8'b10110100} :
//               (x1 == 4'b1111 && x2 == 4'b1101) ? {8'b11000011} :
//               (x1 == 4'b1111 && x2 == 4'b1110) ? {8'b11010010} : {8'b11100001};
// endmodule

// module mul8
//    (  input wire [7:0]  x1,
//       input wire [7:0]  x2,
//       output wire [15:0] y);
   
//    wire [7:0] y1;
//    wire [7:0] y21;
//    wire [7:0] y22;
//    wire [7:0] y3;
//    mul4 u1(x1[3:0],x2[3:0],y1);
//    mul4 u2(x1[3:0],x2[7:4],y21);
//    mul4 u3(x1[7:4],x2[3:0],y22);
//    mul4 u4(x1[7:4],x2[7:4],y3);
//    assign y = {y3,8'b0} + {4'b0,y21,4'b0} + {4'b0,y22,4'b0} + {8'b0,y1};
// endmodule

// module mul16
//    (  input wire [15:0]  x1,
//       input wire [15:0]  x2,
//       output wire [31:0] y);
   
//    wire [15:0] y1;
//    wire [15:0] y21;
//    wire [15:0] y22;
//    wire [15:0] y3;
//    mul8 u1(x1[7:0],x2[7:0],y1);
//    mul8 u2(x1[7:0],x2[15:8],y21);
//    mul8 u3(x1[15:8],x2[7:0],y22);
//    mul8 u4(x1[15:8],x2[15:8],y3);
//    assign y = {y3,16'b0} + {8'b0,y21,8'b0} + {8'b0,y22,8'b0} + {16'b0,y1};
// endmodule

module mul
   (  input wire [31:0]  x1,
      input wire [31:0]  x2,
      output wire [31:0] y,
      output wire        ovf);
   
   // wire [31:0] y1;
   // wire [31:0] y21;
   // wire [31:0] y22;
   // mul16 u1(x1[15:0],x2[15:0],y1);
   // mul16 u2(x1[15:0],x2[31:16],y21);
   // mul16 u3(x1[31:16],x2[15:0],y22);
   // // y1 の32桁目，y21, y22 の 16桁目の内少なくとも2つは0のとき
   // wire [32:0] yl = {y21[15:0],16'b0} + {y22[15:0],16'b0} + y1;

   wire [31:0] y1 = x1[15:0] * x2[15:0];
   wire [31:0] y21 = x1[15:0] * x2[31:16];
   wire [31:0] y22 = x1[31:16] * x2[15:0];
   wire [32:0] yl = {y21[15:0],16'b0} + {y22[15:0],16'b0} + y1;

   assign y = yl[31:0];

   assign ovf = ((|x1[31:16] && |x2[31:16]) || (y1[31:31] && y21[15:15]) || (y1[31:31] && y22[15:15]) || (y21[15:15] && y22[15:15]) || yl[32:32]) ? 1'b1 : 1'b0;

endmodule                                                                         
`default_nettype wire