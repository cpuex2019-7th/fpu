`default_nettype none

module finv
   (  input wire [31:0]  x,
      output wire [31:0] y,
      output wire        exception);
   // 定義
   wire s = x[31:31];
   wire [7:0] e = x[30:23];
   // wire [22:0] m = x[22:0];
   // 非正規化数はinfになるので無視 小数点以下23桁
   wire [23:0] ma = {1'b1,x[22:0]};
   assign [7:0] e3 = e;
   assign s3 = s;
   assign [23:0] ma1 = ma;
   assign [31:0] x3 = x;

   // 小数点以下26
   wire [25:0] x_in = (ma1[22:15] == 8'b00000000) ? {26'b11111111100000000011111111} :
                      (ma1[22:15] == 8'b00000001) ? {26'b11111110100000100011110010} :
                      (ma1[22:15] == 8'b00000010) ? {26'b11111101100001100011000010} :
                      (ma1[22:15] == 8'b00000011) ? {26'b11111100100011000001010110} :
                      (ma1[22:15] == 8'b00000100) ? {26'b11111011100100111110011001} :
                      (ma1[22:15] == 8'b00000101) ? {26'b11111010100111011001110100} :
                      (ma1[22:15] == 8'b00000110) ? {26'b11111001101010010011010000} :
                      (ma1[22:15] == 8'b00000111) ? {26'b11111000101101101010011000} :
                      (ma1[22:15] == 8'b00001000) ? {26'b11110111110001011110110110} :
                      (ma1[22:15] == 8'b00001001) ? {26'b11110110110101110000010101} :
                      (ma1[22:15] == 8'b00001010) ? {26'b11110101111010011110011111} :
                      (ma1[22:15] == 8'b00001011) ? {26'b11110100111111101001000010} :
                      (ma1[22:15] == 8'b00001100) ? {26'b11110100000101001111100111} :
                      (ma1[22:15] == 8'b00001101) ? {26'b11110011001011010001111011} :
                      (ma1[22:15] == 8'b00001110) ? {26'b11110010010001101111101011} :
                      (ma1[22:15] == 8'b00001111) ? {26'b11110001011000101000100010} :
                      (ma1[22:15] == 8'b00010000) ? {26'b11110000011111111100001111} :
                      (ma1[22:15] == 8'b00010001) ? {26'b11101111100111101010011110} :
                      (ma1[22:15] == 8'b00010010) ? {26'b11101110101111110010111100} :
                      (ma1[22:15] == 8'b00010011) ? {26'b11101101111000010101010111} :
                      (ma1[22:15] == 8'b00010100) ? {26'b11101101000001010001011110} :
                      (ma1[22:15] == 8'b00010101) ? {26'b11101100001010100110111110} :
                      (ma1[22:15] == 8'b00010110) ? {26'b11101011010100010101100110} :
                      (ma1[22:15] == 8'b00010111) ? {26'b11101010011110011101000101} :
                      (ma1[22:15] == 8'b00011000) ? {26'b11101001101000111101001001} :
                      (ma1[22:15] == 8'b00011001) ? {26'b11101000110011110101100010} :
                      (ma1[22:15] == 8'b00011010) ? {26'b11100111111111000110000000} :
                      (ma1[22:15] == 8'b00011011) ? {26'b11100111001010101110010001} :
                      (ma1[22:15] == 8'b00011100) ? {26'b11100110010110101110000111} :
                      (ma1[22:15] == 8'b00011101) ? {26'b11100101100011000101010001} :
                      (ma1[22:15] == 8'b00011110) ? {26'b11100100101111110011011111} :
                      (ma1[22:15] == 8'b00011111) ? {26'b11100011111100111000100010} :
                      (ma1[22:15] == 8'b00100000) ? {26'b11100011001010010100001011} :
                      (ma1[22:15] == 8'b00100001) ? {26'b11100010011000000110001100} :
                      (ma1[22:15] == 8'b00100010) ? {26'b11100001100110001110010100} :
                      (ma1[22:15] == 8'b00100011) ? {26'b11100000110100101100010110} :
                      (ma1[22:15] == 8'b00100100) ? {26'b11100000000011100000000011} :
                      (ma1[22:15] == 8'b00100101) ? {26'b11011111010010101001001101} :
                      (ma1[22:15] == 8'b00100110) ? {26'b11011110100010000111100110} :
                      (ma1[22:15] == 8'b00100111) ? {26'b11011101110001111011000001} :
                      (ma1[22:15] == 8'b00101000) ? {26'b11011101000010000011001111} :
                      (ma1[22:15] == 8'b00101001) ? {26'b11011100010010100000000011} :
                      (ma1[22:15] == 8'b00101010) ? {26'b11011011100011010001010000} :
                      (ma1[22:15] == 8'b00101011) ? {26'b11011010110100010110101001} :
                      (ma1[22:15] == 8'b00101100) ? {26'b11011010000101110000000001} :
                      (ma1[22:15] == 8'b00101101) ? {26'b11011001010111011101001011} :
                      (ma1[22:15] == 8'b00101110) ? {26'b11011000101001011101111011} :
                      (ma1[22:15] == 8'b00101111) ? {26'b11010111111011110010000101} :
                      (ma1[22:15] == 8'b00110000) ? {26'b11010111001110011001011011} :
                      (ma1[22:15] == 8'b00110001) ? {26'b11010110100001010011110011} :
                      (ma1[22:15] == 8'b00110010) ? {26'b11010101110100100000111111} :
                      (ma1[22:15] == 8'b00110011) ? {26'b11010101001000000000110101} :
                      (ma1[22:15] == 8'b00110100) ? {26'b11010100011011110011001000} :
                      (ma1[22:15] == 8'b00110101) ? {26'b11010011101111110111101110} :
                      (ma1[22:15] == 8'b00110110) ? {26'b11010011000100001110011011} :
                      (ma1[22:15] == 8'b00110111) ? {26'b11010010011000110111000100} :
                      (ma1[22:15] == 8'b00111000) ? {26'b11010001101101110001011101} :
                      (ma1[22:15] == 8'b00111001) ? {26'b11010001000010111101011100} :
                      (ma1[22:15] == 8'b00111010) ? {26'b11010000011000011010110111} :
                      (ma1[22:15] == 8'b00111011) ? {26'b11001111101110001001100010} :
                      (ma1[22:15] == 8'b00111100) ? {26'b11001111000100001001010011} :
                      (ma1[22:15] == 8'b00111101) ? {26'b11001110011010011010000000} :
                      (ma1[22:15] == 8'b00111110) ? {26'b11001101110000111011011110} :
                      (ma1[22:15] == 8'b00111111) ? {26'b11001101000111101101100100} :
                      (ma1[22:15] == 8'b01000000) ? {26'b11001100011110110000000111} :
                      (ma1[22:15] == 8'b01000001) ? {26'b11001011110110000010111111} :
                      (ma1[22:15] == 8'b01000010) ? {26'b11001011001101100110000000} :
                      (ma1[22:15] == 8'b01000011) ? {26'b11001010100101011001000001} :
                      (ma1[22:15] == 8'b01000100) ? {26'b11001001111101011011111010} :
                      (ma1[22:15] == 8'b01000101) ? {26'b11001001010101101110100000} :
                      (ma1[22:15] == 8'b01000110) ? {26'b11001000101110010000101010} :
                      (ma1[22:15] == 8'b01000111) ? {26'b11001000000111000010001111} :
                      (ma1[22:15] == 8'b01001000) ? {26'b11000111100000000011000111} :
                      (ma1[22:15] == 8'b01001001) ? {26'b11000110111001010011001000} :
                      (ma1[22:15] == 8'b01001010) ? {26'b11000110010010110010001001} :
                      (ma1[22:15] == 8'b01001011) ? {26'b11000101101100100000000011} :
                      (ma1[22:15] == 8'b01001100) ? {26'b11000101000110011100101011} :
                      (ma1[22:15] == 8'b01001101) ? {26'b11000100100000100111111010} :
                      (ma1[22:15] == 8'b01001110) ? {26'b11000011111011000001101000} :
                      (ma1[22:15] == 8'b01001111) ? {26'b11000011010101101001101011} :
                      (ma1[22:15] == 8'b01010000) ? {26'b11000010110000011111111100} :
                      (ma1[22:15] == 8'b01010001) ? {26'b11000010001011100100010100} :
                      (ma1[22:15] == 8'b01010010) ? {26'b11000001100110110110101001} :
                      (ma1[22:15] == 8'b01010011) ? {26'b11000001000010010110110011} :
                      (ma1[22:15] == 8'b01010100) ? {26'b11000000011110000100101100} :
                      (ma1[22:15] == 8'b01010101) ? {26'b10111111111010000000001011} :
                      (ma1[22:15] == 8'b01010110) ? {26'b10111111010110001001001001} :
                      (ma1[22:15] == 8'b01010111) ? {26'b10111110110010011111011111} :
                      (ma1[22:15] == 8'b01011000) ? {26'b10111110001111000011000100} :
                      (ma1[22:15] == 8'b01011001) ? {26'b10111101101011110011110001} :
                      (ma1[22:15] == 8'b01011010) ? {26'b10111101001000110001100000} :
                      (ma1[22:15] == 8'b01011011) ? {26'b10111100100101111100001000} :
                      (ma1[22:15] == 8'b01011100) ? {26'b10111100000011010011100011} :
                      (ma1[22:15] == 8'b01011101) ? {26'b10111011100000110111101010} :
                      (ma1[22:15] == 8'b01011110) ? {26'b10111010111110101000010110} :
                      (ma1[22:15] == 8'b01011111) ? {26'b10111010011100100101100000} :
                      (ma1[22:15] == 8'b01100000) ? {26'b10111001111010101111000001} :
                      (ma1[22:15] == 8'b01100001) ? {26'b10111001011001000100110011} :
                      (ma1[22:15] == 8'b01100010) ? {26'b10111000110111100110101110} :
                      (ma1[22:15] == 8'b01100011) ? {26'b10111000010110010100101101} :
                      (ma1[22:15] == 8'b01100100) ? {26'b10110111110101001110101000} :
                      (ma1[22:15] == 8'b01100101) ? {26'b10110111010100010100011010} :
                      (ma1[22:15] == 8'b01100110) ? {26'b10110110110011100101111011} :
                      (ma1[22:15] == 8'b01100111) ? {26'b10110110010011000011000111} :
                      (ma1[22:15] == 8'b01101000) ? {26'b10110101110010101011110110} :
                      (ma1[22:15] == 8'b01101001) ? {26'b10110101010010100000000010} :
                      (ma1[22:15] == 8'b01101010) ? {26'b10110100110010011111100110} :
                      (ma1[22:15] == 8'b01101011) ? {26'b10110100010010101010011011} :
                      (ma1[22:15] == 8'b01101100) ? {26'b10110011110011000000011100} :
                      (ma1[22:15] == 8'b01101101) ? {26'b10110011010011100001100010} :
                      (ma1[22:15] == 8'b01101110) ? {26'b10110010110100001101100111} :
                      (ma1[22:15] == 8'b01101111) ? {26'b10110010010101000100100111} :
                      (ma1[22:15] == 8'b01110000) ? {26'b10110001110110000110011011} :
                      (ma1[22:15] == 8'b01110001) ? {26'b10110001010111010010111101} :
                      (ma1[22:15] == 8'b01110010) ? {26'b10110000111000101010001001} :
                      (ma1[22:15] == 8'b01110011) ? {26'b10110000011010001011111000} :
                      (ma1[22:15] == 8'b01110100) ? {26'b10101111111011111000000110} :
                      (ma1[22:15] == 8'b01110101) ? {26'b10101111011101101110101100} :
                      (ma1[22:15] == 8'b01110110) ? {26'b10101110111111101111100110} :
                      (ma1[22:15] == 8'b01110111) ? {26'b10101110100001111010101101} :
                      (ma1[22:15] == 8'b01111000) ? {26'b10101110000100001111111110} :
                      (ma1[22:15] == 8'b01111001) ? {26'b10101101100110101111010011} :
                      (ma1[22:15] == 8'b01111010) ? {26'b10101101001001011000100110} :
                      (ma1[22:15] == 8'b01111011) ? {26'b10101100101100001011110011} :
                      (ma1[22:15] == 8'b01111100) ? {26'b10101100001111001000110101} :
                      (ma1[22:15] == 8'b01111101) ? {26'b10101011110010001111100110} :
                      (ma1[22:15] == 8'b01111110) ? {26'b10101011010101100000000010} :
                      (ma1[22:15] == 8'b01111111) ? {26'b10101010111000111010000100} :
                      (ma1[22:15] == 8'b10000000) ? {26'b10101010011100011101101000} :
                      (ma1[22:15] == 8'b10000001) ? {26'b10101010000000001010101000} :
                      (ma1[22:15] == 8'b10000010) ? {26'b10101001100100000000111111} :
                      (ma1[22:15] == 8'b10000011) ? {26'b10101001001000000000101010} :
                      (ma1[22:15] == 8'b10000100) ? {26'b10101000101100001001100011} :
                      (ma1[22:15] == 8'b10000101) ? {26'b10101000010000011011100110} :
                      (ma1[22:15] == 8'b10000110) ? {26'b10100111110100110110101111} :
                      (ma1[22:15] == 8'b10000111) ? {26'b10100111011001011010111001} :
                      (ma1[22:15] == 8'b10001000) ? {26'b10100110111110000111111111} :
                      (ma1[22:15] == 8'b10001001) ? {26'b10100110100010111101111101} :
                      (ma1[22:15] == 8'b10001010) ? {26'b10100110000111111100110000} :
                      (ma1[22:15] == 8'b10001011) ? {26'b10100101101101000100010010} :
                      (ma1[22:15] == 8'b10001100) ? {26'b10100101010010010100011111} :
                      (ma1[22:15] == 8'b10001101) ? {26'b10100100110111101101010100} :
                      (ma1[22:15] == 8'b10001110) ? {26'b10100100011101001110101100} :
                      (ma1[22:15] == 8'b10001111) ? {26'b10100100000010111000100011} :
                      (ma1[22:15] == 8'b10010000) ? {26'b10100011101000101010110100} :
                      (ma1[22:15] == 8'b10010001) ? {26'b10100011001110100101011101} :
                      (ma1[22:15] == 8'b10010010) ? {26'b10100010110100101000011000} :
                      (ma1[22:15] == 8'b10010011) ? {26'b10100010011010110011100011} :
                      (ma1[22:15] == 8'b10010100) ? {26'b10100010000001000110111000} :
                      (ma1[22:15] == 8'b10010101) ? {26'b10100001100111100010010100} :
                      (ma1[22:15] == 8'b10010110) ? {26'b10100001001110000101110100} :
                      (ma1[22:15] == 8'b10010111) ? {26'b10100000110100110001010100} :
                      (ma1[22:15] == 8'b10011000) ? {26'b10100000011011100100101111} :
                      (ma1[22:15] == 8'b10011001) ? {26'b10100000000010100000000010} :
                      (ma1[22:15] == 8'b10011010) ? {26'b10011111101001100011001010} :
                      (ma1[22:15] == 8'b10011011) ? {26'b10011111010000101110000010} :
                      (ma1[22:15] == 8'b10011100) ? {26'b10011110111000000000100111} :
                      (ma1[22:15] == 8'b10011101) ? {26'b10011110011111011010110110} :
                      (ma1[22:15] == 8'b10011110) ? {26'b10011110000110111100101011} :
                      (ma1[22:15] == 8'b10011111) ? {26'b10011101101110100110000010} :
                      (ma1[22:15] == 8'b10100000) ? {26'b10011101010110010110111001} :
                      (ma1[22:15] == 8'b10100001) ? {26'b10011100111110001111001011} :
                      (ma1[22:15] == 8'b10100010) ? {26'b10011100100110001110110101} :
                      (ma1[22:15] == 8'b10100011) ? {26'b10011100001110010101110100} :
                      (ma1[22:15] == 8'b10100100) ? {26'b10011011110110100100000100} :
                      (ma1[22:15] == 8'b10100101) ? {26'b10011011011110111001100010} :
                      (ma1[22:15] == 8'b10100110) ? {26'b10011011000111010110001100} :
                      (ma1[22:15] == 8'b10100111) ? {26'b10011010101111111001111101} :
                      (ma1[22:15] == 8'b10101000) ? {26'b10011010011000100100110010} :
                      (ma1[22:15] == 8'b10101001) ? {26'b10011010000001010110101000} :
                      (ma1[22:15] == 8'b10101010) ? {26'b10011001101010001111011101} :
                      (ma1[22:15] == 8'b10101011) ? {26'b10011001010011001111001100} :
                      (ma1[22:15] == 8'b10101100) ? {26'b10011000111100010101110011} :
                      (ma1[22:15] == 8'b10101101) ? {26'b10011000100101100011001111} :
                      (ma1[22:15] == 8'b10101110) ? {26'b10011000001110110111011100} :
                      (ma1[22:15] == 8'b10101111) ? {26'b10010111111000010010011001} :
                      (ma1[22:15] == 8'b10110000) ? {26'b10010111100001110100000000} :
                      (ma1[22:15] == 8'b10110001) ? {26'b10010111001011011100010001} :
                      (ma1[22:15] == 8'b10110010) ? {26'b10010110110101001011000111} :
                      (ma1[22:15] == 8'b10110011) ? {26'b10010110011111000000100000} :
                      (ma1[22:15] == 8'b10110100) ? {26'b10010110001000111100011010} :
                      (ma1[22:15] == 8'b10110101) ? {26'b10010101110010111110110000} :
                      (ma1[22:15] == 8'b10110110) ? {26'b10010101011101000111100001} :
                      (ma1[22:15] == 8'b10110111) ? {26'b10010101000111010110101001} :
                      (ma1[22:15] == 8'b10111000) ? {26'b10010100110001101100000110} :
                      (ma1[22:15] == 8'b10111001) ? {26'b10010100011100000111110100} :
                      (ma1[22:15] == 8'b10111010) ? {26'b10010100000110101001110011} :
                      (ma1[22:15] == 8'b10111011) ? {26'b10010011110001010001111101} :
                      (ma1[22:15] == 8'b10111100) ? {26'b10010011011100000000010010} :
                      (ma1[22:15] == 8'b10111101) ? {26'b10010011000110110100101110} :
                      (ma1[22:15] == 8'b10111110) ? {26'b10010010110001101111001110} :
                      (ma1[22:15] == 8'b10111111) ? {26'b10010010011100101111110001} :
                      (ma1[22:15] == 8'b11000000) ? {26'b10010010000111110110010010} :
                      (ma1[22:15] == 8'b11000001) ? {26'b10010001110011000010110001} :
                      (ma1[22:15] == 8'b11000010) ? {26'b10010001011110010101001010} :
                      (ma1[22:15] == 8'b11000011) ? {26'b10010001001001101101011011} :
                      (ma1[22:15] == 8'b11000100) ? {26'b10010000110101001011100001} :
                      (ma1[22:15] == 8'b11000101) ? {26'b10010000100000101111011010} :
                      (ma1[22:15] == 8'b11000110) ? {26'b10010000001100011001000100} :
                      (ma1[22:15] == 8'b11000111) ? {26'b10001111111000001000011011} :
                      (ma1[22:15] == 8'b11001000) ? {26'b10001111100011111101011110} :
                      (ma1[22:15] == 8'b11001001) ? {26'b10001111001111111000001010} :
                      (ma1[22:15] == 8'b11001010) ? {26'b10001110111011111000011101} :
                      (ma1[22:15] == 8'b11001011) ? {26'b10001110100111111110010101} :
                      (ma1[22:15] == 8'b11001100) ? {26'b10001110010100001001101110} :
                      (ma1[22:15] == 8'b11001101) ? {26'b10001110000000011010101000} :
                      (ma1[22:15] == 8'b11001110) ? {26'b10001101101100110000111111} :
                      (ma1[22:15] == 8'b11001111) ? {26'b10001101011001001100110001} :
                      (ma1[22:15] == 8'b11010000) ? {26'b10001101000101101101111100} :
                      (ma1[22:15] == 8'b11010001) ? {26'b10001100110010010100011111} :
                      (ma1[22:15] == 8'b11010010) ? {26'b10001100011111000000010101} :
                      (ma1[22:15] == 8'b11010011) ? {26'b10001100001011110001011111} :
                      (ma1[22:15] == 8'b11010100) ? {26'b10001011111000100111111000} :
                      (ma1[22:15] == 8'b11010101) ? {26'b10001011100101100011100000} :
                      (ma1[22:15] == 8'b11010110) ? {26'b10001011010010100100010100} :
                      (ma1[22:15] == 8'b11010111) ? {26'b10001010111111101010010010} :
                      (ma1[22:15] == 8'b11011000) ? {26'b10001010101100110101010111} :
                      (ma1[22:15] == 8'b11011001) ? {26'b10001010011010000101100010} :
                      (ma1[22:15] == 8'b11011010) ? {26'b10001010000111011010110001} :
                      (ma1[22:15] == 8'b11011011) ? {26'b10001001110100110101000001} :
                      (ma1[22:15] == 8'b11011100) ? {26'b10001001100010010100010001} :
                      (ma1[22:15] == 8'b11011101) ? {26'b10001001001111111000011111} :
                      (ma1[22:15] == 8'b11011110) ? {26'b10001000111101100001101000} :
                      (ma1[22:15] == 8'b11011111) ? {26'b10001000101011001111101011} :
                      (ma1[22:15] == 8'b11100000) ? {26'b10001000011001000010100110} :
                      (ma1[22:15] == 8'b11100001) ? {26'b10001000000110111010010110} :
                      (ma1[22:15] == 8'b11100010) ? {26'b10000111110100110110111010} :
                      (ma1[22:15] == 8'b11100011) ? {26'b10000111100010111000010000} :
                      (ma1[22:15] == 8'b11100100) ? {26'b10000111010000111110010110} :
                      (ma1[22:15] == 8'b11100101) ? {26'b10000110111111001001001010} :
                      (ma1[22:15] == 8'b11100110) ? {26'b10000110101101011000101010} :
                      (ma1[22:15] == 8'b11100111) ? {26'b10000110011011101100110101} :
                      (ma1[22:15] == 8'b11101000) ? {26'b10000110001010000101101000} :
                      (ma1[22:15] == 8'b11101001) ? {26'b10000101111000100011000010} :
                      (ma1[22:15] == 8'b11101010) ? {26'b10000101100111000101000001} :
                      (ma1[22:15] == 8'b11101011) ? {26'b10000101010101101011100011} :
                      (ma1[22:15] == 8'b11101100) ? {26'b10000101000100010110100111} :
                      (ma1[22:15] == 8'b11101101) ? {26'b10000100110011000110001010} :
                      (ma1[22:15] == 8'b11101110) ? {26'b10000100100001111010001011} :
                      (ma1[22:15] == 8'b11101111) ? {26'b10000100010000110010101000} :
                      (ma1[22:15] == 8'b11110000) ? {26'b10000011111111101111100000} :
                      (ma1[22:15] == 8'b11110001) ? {26'b10000011101110110000110000} :
                      (ma1[22:15] == 8'b11110010) ? {26'b10000011011101110110010111} :
                      (ma1[22:15] == 8'b11110011) ? {26'b10000011001101000000010100} :
                      (ma1[22:15] == 8'b11110100) ? {26'b10000010111100001110100100} :
                      (ma1[22:15] == 8'b11110101) ? {26'b10000010101011100001000111} :
                      (ma1[22:15] == 8'b11110110) ? {26'b10000010011010110111111010} :
                      (ma1[22:15] == 8'b11110111) ? {26'b10000010001010010010111100} :
                      (ma1[22:15] == 8'b11111000) ? {26'b10000001111001110010001011} :
                      (ma1[22:15] == 8'b11111001) ? {26'b10000001101001010101100101} :
                      (ma1[22:15] == 8'b11111010) ? {26'b10000001011000111101001010} :
                      (ma1[22:15] == 8'b11111011) ? {26'b10000001001000101000110110} :
                      (ma1[22:15] == 8'b11111100) ? {26'b10000000111000011000101010} :
                      (ma1[22:15] == 8'b11111101) ? {26'b10000000101000001100100011} :
                      (ma1[22:15] == 8'b11111110) ? {26'b10000000011000000100100000} : {26'b10000000001000000000100000};

   // ニュートン法1回目
   // x_out1 = x_in*(2-a*x_in)
   // x_in*(2-a*x_in) 小数点以下75桁
   wire [74:0] k1 = {51'b0,ma1} * {49'b0,x_in} * {49'b0,x_in};
   wire [75:0] p1 = {x_in,50'b0} - {1'b0,k1};
   // 切り上げるのは p1[48]が1かつ(p1[47:0]が0より大きい または p1[49]が1)
   // 上二桁が整数部
   wire [25:0] x_out1 = (p1[48:48] && (|p1[47:0] || p1[49:49])) ? {p1[74:49]} + 26'b1 : {p1[74:49]};
   assign [25:0] x_out11 = x_out1;
   assign [7:0] e4 = e;
   assign s4 = s;
   assign [23:0] ma2 = ma;
   assign [31:0] x4 = x;

   // ニュートン法2回目
   wire [74:0] k2 = {51'b0,ma2} * {49'b0,x_out11} * {49'b0,x_out11};
   wire [75:0] p2 = {x_out11,50'b0} - {1'b0,k2};
   wire [25:0] x_out2 = (p2[48:48] && (|p2[47:0] || p2[49:49])) ? {p2[74:49]} + 26'b1 : {p2[74:49]};

   wire [22:0] my = (e4 == 8'd254) ? ((x_out2[3:3]) ? {1'b0,x_out2[25:4]} + 23'b1 : {1'b0,x_out2[25:4]}) :
                    (e4 == 8'd253) ? ((x_out2[2:2]) ? x_out2[25:3] + 23'b1 : x_out2[25:3]) :
                    (x_out2[1:1]) ? x_out2[24:2] + 23'b1 : x_out2[24:2];

   wire [7:0] ey = (e4 == 8'd254) ? 0 : 8'd253 - e4;
   wire [7:0] ey2 = (e4 == 8'd253) ? 0 : ey + 8'b1;

   // nanかどうかの判定
   wire nzm = |x4[22:0];
   assign y = (e4 == 8'd255 && nzm) ? {s4,8'd255,1'b1,x4[21:0]} : // 元がnanなら結果もnan
              (e4 == 8'd255 && ~nzm) ? {s4,8'd0,23'b0} : // 元がinfなら結果は0
              (~|x4) ? {s4,8'd255,23'b0} : // 元が+-0なら結果は+-inf
              (~|x4[22:0]) ? ((e4 == 8'd254) ? {s4,8'b0,1'b1,22'b0} : (e4 == 8'd253) ? {s4,8'b1,23'b0} : {s4,ey2,23'b0}) : {s4,ey,my};

   assign exception = (e4 == 8'd255 && nzm) ? 1'b1 : 1'b0;

endmodule

module fdiv
   (  input wire [31:0]  x1,
      input wire [31:0]  x2,
      output wire [31:0] y,
      output wire        ovf);
   // 定義
   wire s1 = x1[31:31];
   wire [7:0] e1 = x1[30:23];
   wire [22:0] m1 = x1[22:0];
   wire s2 = x2[31:31];
   wire [7:0] e2 = x2[30:23];
   wire [22:0] m2 = x2[22:0];

   wire [31:0] x2i;
   wire exception;
   finv u1(x2,x2i,exception);
   assign [31:0] y1 = y;
   assign [31:0] x11 = x1;
   fmul u2(x2i,x1,y,ovf);

endmodule                                                                         
`default_nettype wire