`default_nettype none

module fmul
   (  input wire [31:0]  x1,
      input wire [31:0]  x2,
      output wire [31:0] y,
      output wire        ovf);
   // 定義
   wire s1 = x1[31:31];
   wire [7:0] e1 = x1[30:23];
   wire [22:0] m1 = x1[22:0];
   wire s2 = x2[31:31];
   wire [7:0] e2 = x2[30:23];
   wire [22:0] m2 = x2[22:0];
   // 非正規化数の処理
   wire [23:0] m1a = (e1 == 8'b0) ? {1'b0,m1} : {1'b1,m1};
   wire [23:0] m2a = (e2 == 8'b0) ? {1'b0,m2} : {1'b1,m2};
   wire [7:0] e1a = (e1 == 8'b0) ? 8'b1 : e1;
   wire [7:0] e2a = (e2 == 8'b0) ? 8'b1 : e2;
   // mantissaの掛け算の計算
   wire [47:0] mye = {24'b0,m1a} * {24'b0,m2a};
   // 何桁ずらすかを計算
   wire [5:0] se = (mye[47:47]) ? 6'd0 :
                   (mye[46:46]) ? 6'd1 :
                   (mye[45:45]) ? 6'd2 :
                   (mye[44:44]) ? 6'd3 :
                   (mye[43:43]) ? 6'd4 :
                   (mye[42:42]) ? 6'd5 :
                   (mye[41:41]) ? 6'd6 :
                   (mye[40:40]) ? 6'd7 :
                   (mye[39:39]) ? 6'd8 :
                   (mye[38:38]) ? 6'd9 :
                   (mye[37:37]) ? 6'd10 :
                   (mye[36:36]) ? 6'd11 :
                   (mye[35:35]) ? 6'd12 :
                   (mye[34:34]) ? 6'd13 :
                   (mye[33:33]) ? 6'd14 :
                   (mye[32:32]) ? 6'd15 :
                   (mye[31:31]) ? 6'd16 :
                   (mye[30:30]) ? 6'd17 :
                   (mye[29:29]) ? 6'd18 :
                   (mye[28:28]) ? 6'd19 :
                   (mye[27:27]) ? 6'd20 :
                   (mye[26:26]) ? 6'd21 :
                   (mye[25:25]) ? 6'd22 :
                   (mye[24:24]) ? 6'd23 :
                   (mye[23:23]) ? 6'd24 :
                   (mye[22:22]) ? 6'd25 :
                   (mye[21:21]) ? 6'd26 :
                   (mye[20:20]) ? 6'd27 :
                   (mye[19:19]) ? 6'd28 :
                   (mye[18:18]) ? 6'd29 :
                   (mye[17:17]) ? 6'd30 :
                   (mye[16:16]) ? 6'd31 :
                   (mye[15:15]) ? 6'd32 :
                   (mye[14:14]) ? 6'd33 :
                   (mye[13:13]) ? 6'd34 :
                   (mye[12:12]) ? 6'd35 :
                   (mye[11:11]) ? 6'd36 :
                   (mye[10:10]) ? 6'd37 :
                   (mye[9:9]) ? 6'd38 :
                   (mye[8:8]) ? 6'd39 :
                   (mye[7:7]) ? 6'd40 :
                   (mye[6:6]) ? 6'd41 :
                   (mye[5:5]) ? 6'd42 :
                   (mye[4:4]) ? 6'd43 :
                   (mye[3:3]) ? 6'd44 :
                   (mye[2:2]) ? 6'd45 :
                   (mye[1:1]) ? 6'd46 :
                   (mye[0:0]) ? 6'd47 : 6'd48;
   // myft[47]に1が来るように左シフト
   wire [47:0] myft = (mye[47:47]) ? mye :
                      (mye[46:46]) ? {mye[46:0],1'b0} :
                      (mye[45:45]) ? {mye[45:0],2'b0} :
                      (mye[44:44]) ? {mye[44:0],3'b0} :
                      (mye[43:43]) ? {mye[43:0],4'b0} :
                      (mye[42:42]) ? {mye[42:0],5'b0} :
                      (mye[41:41]) ? {mye[41:0],6'b0} :
                      (mye[40:40]) ? {mye[40:0],7'b0} :
                      (mye[39:39]) ? {mye[39:0],8'b0} :
                      (mye[38:38]) ? {mye[38:0],9'b0} :
                      (mye[37:37]) ? {mye[37:0],10'b0} :
                      (mye[36:36]) ? {mye[36:0],11'b0} :
                      (mye[35:35]) ? {mye[35:0],12'b0} :
                      (mye[34:34]) ? {mye[34:0],13'b0} :
                      (mye[33:33]) ? {mye[33:0],14'b0} :
                      (mye[32:32]) ? {mye[32:0],15'b0} :
                      (mye[31:31]) ? {mye[31:0],16'b0} :
                      (mye[30:30]) ? {mye[30:0],17'b0} :
                      (mye[29:29]) ? {mye[29:0],18'b0} :
                      (mye[28:28]) ? {mye[28:0],19'b0} :
                      (mye[27:27]) ? {mye[27:0],20'b0} :
                      (mye[26:26]) ? {mye[26:0],21'b0} :
                      (mye[25:25]) ? {mye[25:0],22'b0} :
                      (mye[24:24]) ? {mye[24:0],23'b0} :
                      (mye[23:23]) ? {mye[23:0],24'b0} :
                      (mye[22:22]) ? {mye[22:0],25'b0} :
                      (mye[21:21]) ? {mye[21:0],26'b0} :
                      (mye[20:20]) ? {mye[20:0],27'b0} :
                      (mye[19:19]) ? {mye[19:0],28'b0} :
                      (mye[18:18]) ? {mye[18:0],29'b0} :
                      (mye[17:17]) ? {mye[17:0],30'b0} :
                      (mye[16:16]) ? {mye[16:0],31'b0} :
                      (mye[15:15]) ? {mye[15:0],32'b0} :
                      (mye[14:14]) ? {mye[14:0],33'b0} :
                      (mye[13:13]) ? {mye[13:0],34'b0} :
                      (mye[12:12]) ? {mye[12:0],35'b0} :
                      (mye[11:11]) ? {mye[11:0],36'b0} :
                      (mye[10:10]) ? {mye[10:0],37'b0} :
                      (mye[9:9]) ? {mye[9:0],38'b0} :
                      (mye[8:8]) ? {mye[8:0],39'b0} :
                      (mye[7:7]) ? {mye[7:0],40'b0} :
                      (mye[6:6]) ? {mye[6:0],41'b0} :
                      (mye[5:5]) ? {mye[5:0],42'b0} :
                      (mye[4:4]) ? {mye[4:0],43'b0} :
                      (mye[3:3]) ? {mye[3:0],44'b0} :
                      (mye[2:2]) ? {mye[2:0],45'b0} :
                      (mye[1:1]) ? {mye[1:0],46'b0} :
                      (mye[0:0]) ? {mye[0:0],47'b0} : 48'b0;
   // seが0のとき1繰り上がり，そうでないときはse-1繰り下がる
   wire [9:0] eyrt = {2'b0,e1a} + {2'b0,e2a} - {4'b0,se} - 10'd126;
   wire [7:0] eyr = (eyrt[9:9]) ? 8'b0 : (eyrt[8:8]) ? 8'd255 : eyrt[7:0];
   // eyri = eyr + 1
   wire [9:0] eyrit = eyrt + 10'b1;
   wire [7:0] eyri = (eyrit[9:9]) ? 8'b0 : (eyrit[8:8]) ? 8'd255 : eyrit[7:0];
   // eyrtが負のとき正規化するためにmyeをss右シフト，その他のときはそのまま
   // myft[69:47]がmantissa，myft[46:0]が切り捨てられる部分
   wire [9:0] ss = ~eyrt + 10'd2;
   wire [70:0] myf = (eyrt[9:9]) ? {myft,23'b0} >> ss[7:0] : (~|eyrt) ? {myft,23'b0} >> 1'b1 : {myft,23'b0};
   
   // 偶数丸めを行う
   // 切り上げるのは myf[46]が1かつ(myf[45:0]が0より大きいとき または myf[47]が1のとき)
   wire [24:0] myr = (myf[46:46]) ? {1'b0,myf[70:47]} + 25'b1 : {1'b0,myf[70:47]};
   // もう一度丸める
   wire [7:0] ey = (myr[24:24] == 1'b1) ? eyri : (myr[23:23] && ~|eyr) ? 8'b1 : (|myr[23:0] == 1'b0) ? 8'b0 : eyr;
   wire [22:0] my = (myr[24:24] == 1'b1) ? 23'b0 : (myr[23:23] && ~|eyr) ? {myr[21:0],1'b0} : myr[22:0];
   // 符号を求める
   wire sy = s1 ^ s2;
   // nanかどうかの判定
   wire nzm1 = |m1;
   wire nzm2 = |m2;
   assign y = (e2 == 8'd255 && nzm2) ? {s2,8'd255,1'b1,m2[21:0]} :
              (e1 == 8'd255 && nzm1) ? {s1,8'd255,1'b1,m1[21:0]} : // 片方がnanなら結果もnan
              (e1 == 8'd255 && e2 == 8'd0 && ~nzm2) ? {1'b1,8'd255,1'b1,m1[21:0]} :
              (e2 == 8'd255 && e1 == 8'd0 && ~nzm1) ? {1'b1,8'd255,1'b1,m2[21:0]} : // 0*infなら-nan
              (e1 == 8'd255 || e2 == 8'd255) ? {sy,8'd255,23'b0} : // 両方無限なら符号を合わせて無限にする
              (e1 < 8'd255 && e2 < 8'd255 && ey == 8'd255) ? {sy,8'd255,23'b0} : {sy,ey,my}; // overflowしたら符号を合わせて無限にする
   assign ovf = (e1 < 8'd255 && e2 < 8'd255 && ey == 8'd255) ? 1'b1 : 1'b0;

endmodule                      

module newton_inv
   ( input wire [23:0] a,
     input wire [25:0] x_in,
     output wire [25:0] x_out);

   // x_out = x_in*(2-a*x_in)
   // x_in*(2-a*x_in) 小数点以下75桁
   wire [74:0] k = {51'b0,a} * {49'b0,x_in} * {49'b0,x_in};
   wire [75:0] p = {x_in,50'b0} - {1'b0,k};

   // 切り上げるのは p[48]が1かつ(p[47:0]が0より大きい または p[49]が1)
   // 上二桁が整数部
   assign x_out = (p[48:48] && (|p[47:0] || p[49:49])) ? {p[74:49]} + 26'b1 : {p[74:49]};

endmodule

module finv
   (  input wire [31:0]  x,
      output wire [31:0] y,
      output wire        exception);
   // 定義
   wire s = x[31:31];
   wire [7:0] e = x[30:23];
   // wire [22:0] m = x[22:0];
   // 非正規化数はinfになるので無視 小数点以下23桁
   wire [23:0] ma = {1'b1,x[22:0]};

   // 小数点以下26
   wire [25:0] x_out0 = (ma[22:15] == 8'b00000000) ? {26'b11111111100000000011111111} :
                        (ma[22:15] == 8'b00000001) ? {26'b11111110100000100011110010} :
                        (ma[22:15] == 8'b00000010) ? {26'b11111101100001100011000010} :
                        (ma[22:15] == 8'b00000011) ? {26'b11111100100011000001010110} :
                        (ma[22:15] == 8'b00000100) ? {26'b11111011100100111110011001} :
                        (ma[22:15] == 8'b00000101) ? {26'b11111010100111011001110100} :
                        (ma[22:15] == 8'b00000110) ? {26'b11111001101010010011010000} :
                        (ma[22:15] == 8'b00000111) ? {26'b11111000101101101010011000} :
                        (ma[22:15] == 8'b00001000) ? {26'b11110111110001011110110110} :
                        (ma[22:15] == 8'b00001001) ? {26'b11110110110101110000010101} :
                        (ma[22:15] == 8'b00001010) ? {26'b11110101111010011110011111} :
                        (ma[22:15] == 8'b00001011) ? {26'b11110100111111101001000010} :
                        (ma[22:15] == 8'b00001100) ? {26'b11110100000101001111100111} :
                        (ma[22:15] == 8'b00001101) ? {26'b11110011001011010001111011} :
                        (ma[22:15] == 8'b00001110) ? {26'b11110010010001101111101011} :
                        (ma[22:15] == 8'b00001111) ? {26'b11110001011000101000100010} :
                        (ma[22:15] == 8'b00010000) ? {26'b11110000011111111100001111} :
                        (ma[22:15] == 8'b00010001) ? {26'b11101111100111101010011110} :
                        (ma[22:15] == 8'b00010010) ? {26'b11101110101111110010111100} :
                        (ma[22:15] == 8'b00010011) ? {26'b11101101111000010101010111} :
                        (ma[22:15] == 8'b00010100) ? {26'b11101101000001010001011110} :
                        (ma[22:15] == 8'b00010101) ? {26'b11101100001010100110111110} :
                        (ma[22:15] == 8'b00010110) ? {26'b11101011010100010101100110} :
                        (ma[22:15] == 8'b00010111) ? {26'b11101010011110011101000101} :
                        (ma[22:15] == 8'b00011000) ? {26'b11101001101000111101001001} :
                        (ma[22:15] == 8'b00011001) ? {26'b11101000110011110101100010} :
                        (ma[22:15] == 8'b00011010) ? {26'b11100111111111000110000000} :
                        (ma[22:15] == 8'b00011011) ? {26'b11100111001010101110010001} :
                        (ma[22:15] == 8'b00011100) ? {26'b11100110010110101110000111} :
                        (ma[22:15] == 8'b00011101) ? {26'b11100101100011000101010001} :
                        (ma[22:15] == 8'b00011110) ? {26'b11100100101111110011011111} :
                        (ma[22:15] == 8'b00011111) ? {26'b11100011111100111000100010} :
                        (ma[22:15] == 8'b00100000) ? {26'b11100011001010010100001011} :
                        (ma[22:15] == 8'b00100001) ? {26'b11100010011000000110001100} :
                        (ma[22:15] == 8'b00100010) ? {26'b11100001100110001110010100} :
                        (ma[22:15] == 8'b00100011) ? {26'b11100000110100101100010110} :
                        (ma[22:15] == 8'b00100100) ? {26'b11100000000011100000000011} :
                        (ma[22:15] == 8'b00100101) ? {26'b11011111010010101001001101} :
                        (ma[22:15] == 8'b00100110) ? {26'b11011110100010000111100110} :
                        (ma[22:15] == 8'b00100111) ? {26'b11011101110001111011000001} :
                        (ma[22:15] == 8'b00101000) ? {26'b11011101000010000011001111} :
                        (ma[22:15] == 8'b00101001) ? {26'b11011100010010100000000011} :
                        (ma[22:15] == 8'b00101010) ? {26'b11011011100011010001010000} :
                        (ma[22:15] == 8'b00101011) ? {26'b11011010110100010110101001} :
                        (ma[22:15] == 8'b00101100) ? {26'b11011010000101110000000001} :
                        (ma[22:15] == 8'b00101101) ? {26'b11011001010111011101001011} :
                        (ma[22:15] == 8'b00101110) ? {26'b11011000101001011101111011} :
                        (ma[22:15] == 8'b00101111) ? {26'b11010111111011110010000101} :
                        (ma[22:15] == 8'b00110000) ? {26'b11010111001110011001011011} :
                        (ma[22:15] == 8'b00110001) ? {26'b11010110100001010011110011} :
                        (ma[22:15] == 8'b00110010) ? {26'b11010101110100100000111111} :
                        (ma[22:15] == 8'b00110011) ? {26'b11010101001000000000110101} :
                        (ma[22:15] == 8'b00110100) ? {26'b11010100011011110011001000} :
                        (ma[22:15] == 8'b00110101) ? {26'b11010011101111110111101110} :
                        (ma[22:15] == 8'b00110110) ? {26'b11010011000100001110011011} :
                        (ma[22:15] == 8'b00110111) ? {26'b11010010011000110111000100} :
                        (ma[22:15] == 8'b00111000) ? {26'b11010001101101110001011101} :
                        (ma[22:15] == 8'b00111001) ? {26'b11010001000010111101011100} :
                        (ma[22:15] == 8'b00111010) ? {26'b11010000011000011010110111} :
                        (ma[22:15] == 8'b00111011) ? {26'b11001111101110001001100010} :
                        (ma[22:15] == 8'b00111100) ? {26'b11001111000100001001010011} :
                        (ma[22:15] == 8'b00111101) ? {26'b11001110011010011010000000} :
                        (ma[22:15] == 8'b00111110) ? {26'b11001101110000111011011110} :
                        (ma[22:15] == 8'b00111111) ? {26'b11001101000111101101100100} :
                        (ma[22:15] == 8'b01000000) ? {26'b11001100011110110000000111} :
                        (ma[22:15] == 8'b01000001) ? {26'b11001011110110000010111111} :
                        (ma[22:15] == 8'b01000010) ? {26'b11001011001101100110000000} :
                        (ma[22:15] == 8'b01000011) ? {26'b11001010100101011001000001} :
                        (ma[22:15] == 8'b01000100) ? {26'b11001001111101011011111010} :
                        (ma[22:15] == 8'b01000101) ? {26'b11001001010101101110100000} :
                        (ma[22:15] == 8'b01000110) ? {26'b11001000101110010000101010} :
                        (ma[22:15] == 8'b01000111) ? {26'b11001000000111000010001111} :
                        (ma[22:15] == 8'b01001000) ? {26'b11000111100000000011000111} :
                        (ma[22:15] == 8'b01001001) ? {26'b11000110111001010011001000} :
                        (ma[22:15] == 8'b01001010) ? {26'b11000110010010110010001001} :
                        (ma[22:15] == 8'b01001011) ? {26'b11000101101100100000000011} :
                        (ma[22:15] == 8'b01001100) ? {26'b11000101000110011100101011} :
                        (ma[22:15] == 8'b01001101) ? {26'b11000100100000100111111010} :
                        (ma[22:15] == 8'b01001110) ? {26'b11000011111011000001101000} :
                        (ma[22:15] == 8'b01001111) ? {26'b11000011010101101001101011} :
                        (ma[22:15] == 8'b01010000) ? {26'b11000010110000011111111100} :
                        (ma[22:15] == 8'b01010001) ? {26'b11000010001011100100010100} :
                        (ma[22:15] == 8'b01010010) ? {26'b11000001100110110110101001} :
                        (ma[22:15] == 8'b01010011) ? {26'b11000001000010010110110011} :
                        (ma[22:15] == 8'b01010100) ? {26'b11000000011110000100101100} :
                        (ma[22:15] == 8'b01010101) ? {26'b10111111111010000000001011} :
                        (ma[22:15] == 8'b01010110) ? {26'b10111111010110001001001001} :
                        (ma[22:15] == 8'b01010111) ? {26'b10111110110010011111011111} :
                        (ma[22:15] == 8'b01011000) ? {26'b10111110001111000011000100} :
                        (ma[22:15] == 8'b01011001) ? {26'b10111101101011110011110001} :
                        (ma[22:15] == 8'b01011010) ? {26'b10111101001000110001100000} :
                        (ma[22:15] == 8'b01011011) ? {26'b10111100100101111100001000} :
                        (ma[22:15] == 8'b01011100) ? {26'b10111100000011010011100011} :
                        (ma[22:15] == 8'b01011101) ? {26'b10111011100000110111101010} :
                        (ma[22:15] == 8'b01011110) ? {26'b10111010111110101000010110} :
                        (ma[22:15] == 8'b01011111) ? {26'b10111010011100100101100000} :
                        (ma[22:15] == 8'b01100000) ? {26'b10111001111010101111000001} :
                        (ma[22:15] == 8'b01100001) ? {26'b10111001011001000100110011} :
                        (ma[22:15] == 8'b01100010) ? {26'b10111000110111100110101110} :
                        (ma[22:15] == 8'b01100011) ? {26'b10111000010110010100101101} :
                        (ma[22:15] == 8'b01100100) ? {26'b10110111110101001110101000} :
                        (ma[22:15] == 8'b01100101) ? {26'b10110111010100010100011010} :
                        (ma[22:15] == 8'b01100110) ? {26'b10110110110011100101111011} :
                        (ma[22:15] == 8'b01100111) ? {26'b10110110010011000011000111} :
                        (ma[22:15] == 8'b01101000) ? {26'b10110101110010101011110110} :
                        (ma[22:15] == 8'b01101001) ? {26'b10110101010010100000000010} :
                        (ma[22:15] == 8'b01101010) ? {26'b10110100110010011111100110} :
                        (ma[22:15] == 8'b01101011) ? {26'b10110100010010101010011011} :
                        (ma[22:15] == 8'b01101100) ? {26'b10110011110011000000011100} :
                        (ma[22:15] == 8'b01101101) ? {26'b10110011010011100001100010} :
                        (ma[22:15] == 8'b01101110) ? {26'b10110010110100001101100111} :
                        (ma[22:15] == 8'b01101111) ? {26'b10110010010101000100100111} :
                        (ma[22:15] == 8'b01110000) ? {26'b10110001110110000110011011} :
                        (ma[22:15] == 8'b01110001) ? {26'b10110001010111010010111101} :
                        (ma[22:15] == 8'b01110010) ? {26'b10110000111000101010001001} :
                        (ma[22:15] == 8'b01110011) ? {26'b10110000011010001011111000} :
                        (ma[22:15] == 8'b01110100) ? {26'b10101111111011111000000110} :
                        (ma[22:15] == 8'b01110101) ? {26'b10101111011101101110101100} :
                        (ma[22:15] == 8'b01110110) ? {26'b10101110111111101111100110} :
                        (ma[22:15] == 8'b01110111) ? {26'b10101110100001111010101101} :
                        (ma[22:15] == 8'b01111000) ? {26'b10101110000100001111111110} :
                        (ma[22:15] == 8'b01111001) ? {26'b10101101100110101111010011} :
                        (ma[22:15] == 8'b01111010) ? {26'b10101101001001011000100110} :
                        (ma[22:15] == 8'b01111011) ? {26'b10101100101100001011110011} :
                        (ma[22:15] == 8'b01111100) ? {26'b10101100001111001000110101} :
                        (ma[22:15] == 8'b01111101) ? {26'b10101011110010001111100110} :
                        (ma[22:15] == 8'b01111110) ? {26'b10101011010101100000000010} :
                        (ma[22:15] == 8'b01111111) ? {26'b10101010111000111010000100} :
                        (ma[22:15] == 8'b10000000) ? {26'b10101010011100011101101000} :
                        (ma[22:15] == 8'b10000001) ? {26'b10101010000000001010101000} :
                        (ma[22:15] == 8'b10000010) ? {26'b10101001100100000000111111} :
                        (ma[22:15] == 8'b10000011) ? {26'b10101001001000000000101010} :
                        (ma[22:15] == 8'b10000100) ? {26'b10101000101100001001100011} :
                        (ma[22:15] == 8'b10000101) ? {26'b10101000010000011011100110} :
                        (ma[22:15] == 8'b10000110) ? {26'b10100111110100110110101111} :
                        (ma[22:15] == 8'b10000111) ? {26'b10100111011001011010111001} :
                        (ma[22:15] == 8'b10001000) ? {26'b10100110111110000111111111} :
                        (ma[22:15] == 8'b10001001) ? {26'b10100110100010111101111101} :
                        (ma[22:15] == 8'b10001010) ? {26'b10100110000111111100110000} :
                        (ma[22:15] == 8'b10001011) ? {26'b10100101101101000100010010} :
                        (ma[22:15] == 8'b10001100) ? {26'b10100101010010010100011111} :
                        (ma[22:15] == 8'b10001101) ? {26'b10100100110111101101010100} :
                        (ma[22:15] == 8'b10001110) ? {26'b10100100011101001110101100} :
                        (ma[22:15] == 8'b10001111) ? {26'b10100100000010111000100011} :
                        (ma[22:15] == 8'b10010000) ? {26'b10100011101000101010110100} :
                        (ma[22:15] == 8'b10010001) ? {26'b10100011001110100101011101} :
                        (ma[22:15] == 8'b10010010) ? {26'b10100010110100101000011000} :
                        (ma[22:15] == 8'b10010011) ? {26'b10100010011010110011100011} :
                        (ma[22:15] == 8'b10010100) ? {26'b10100010000001000110111000} :
                        (ma[22:15] == 8'b10010101) ? {26'b10100001100111100010010100} :
                        (ma[22:15] == 8'b10010110) ? {26'b10100001001110000101110100} :
                        (ma[22:15] == 8'b10010111) ? {26'b10100000110100110001010100} :
                        (ma[22:15] == 8'b10011000) ? {26'b10100000011011100100101111} :
                        (ma[22:15] == 8'b10011001) ? {26'b10100000000010100000000010} :
                        (ma[22:15] == 8'b10011010) ? {26'b10011111101001100011001010} :
                        (ma[22:15] == 8'b10011011) ? {26'b10011111010000101110000010} :
                        (ma[22:15] == 8'b10011100) ? {26'b10011110111000000000100111} :
                        (ma[22:15] == 8'b10011101) ? {26'b10011110011111011010110110} :
                        (ma[22:15] == 8'b10011110) ? {26'b10011110000110111100101011} :
                        (ma[22:15] == 8'b10011111) ? {26'b10011101101110100110000010} :
                        (ma[22:15] == 8'b10100000) ? {26'b10011101010110010110111001} :
                        (ma[22:15] == 8'b10100001) ? {26'b10011100111110001111001011} :
                        (ma[22:15] == 8'b10100010) ? {26'b10011100100110001110110101} :
                        (ma[22:15] == 8'b10100011) ? {26'b10011100001110010101110100} :
                        (ma[22:15] == 8'b10100100) ? {26'b10011011110110100100000100} :
                        (ma[22:15] == 8'b10100101) ? {26'b10011011011110111001100010} :
                        (ma[22:15] == 8'b10100110) ? {26'b10011011000111010110001100} :
                        (ma[22:15] == 8'b10100111) ? {26'b10011010101111111001111101} :
                        (ma[22:15] == 8'b10101000) ? {26'b10011010011000100100110010} :
                        (ma[22:15] == 8'b10101001) ? {26'b10011010000001010110101000} :
                        (ma[22:15] == 8'b10101010) ? {26'b10011001101010001111011101} :
                        (ma[22:15] == 8'b10101011) ? {26'b10011001010011001111001100} :
                        (ma[22:15] == 8'b10101100) ? {26'b10011000111100010101110011} :
                        (ma[22:15] == 8'b10101101) ? {26'b10011000100101100011001111} :
                        (ma[22:15] == 8'b10101110) ? {26'b10011000001110110111011100} :
                        (ma[22:15] == 8'b10101111) ? {26'b10010111111000010010011001} :
                        (ma[22:15] == 8'b10110000) ? {26'b10010111100001110100000000} :
                        (ma[22:15] == 8'b10110001) ? {26'b10010111001011011100010001} :
                        (ma[22:15] == 8'b10110010) ? {26'b10010110110101001011000111} :
                        (ma[22:15] == 8'b10110011) ? {26'b10010110011111000000100000} :
                        (ma[22:15] == 8'b10110100) ? {26'b10010110001000111100011010} :
                        (ma[22:15] == 8'b10110101) ? {26'b10010101110010111110110000} :
                        (ma[22:15] == 8'b10110110) ? {26'b10010101011101000111100001} :
                        (ma[22:15] == 8'b10110111) ? {26'b10010101000111010110101001} :
                        (ma[22:15] == 8'b10111000) ? {26'b10010100110001101100000110} :
                        (ma[22:15] == 8'b10111001) ? {26'b10010100011100000111110100} :
                        (ma[22:15] == 8'b10111010) ? {26'b10010100000110101001110011} :
                        (ma[22:15] == 8'b10111011) ? {26'b10010011110001010001111101} :
                        (ma[22:15] == 8'b10111100) ? {26'b10010011011100000000010010} :
                        (ma[22:15] == 8'b10111101) ? {26'b10010011000110110100101110} :
                        (ma[22:15] == 8'b10111110) ? {26'b10010010110001101111001110} :
                        (ma[22:15] == 8'b10111111) ? {26'b10010010011100101111110001} :
                        (ma[22:15] == 8'b11000000) ? {26'b10010010000111110110010010} :
                        (ma[22:15] == 8'b11000001) ? {26'b10010001110011000010110001} :
                        (ma[22:15] == 8'b11000010) ? {26'b10010001011110010101001010} :
                        (ma[22:15] == 8'b11000011) ? {26'b10010001001001101101011011} :
                        (ma[22:15] == 8'b11000100) ? {26'b10010000110101001011100001} :
                        (ma[22:15] == 8'b11000101) ? {26'b10010000100000101111011010} :
                        (ma[22:15] == 8'b11000110) ? {26'b10010000001100011001000100} :
                        (ma[22:15] == 8'b11000111) ? {26'b10001111111000001000011011} :
                        (ma[22:15] == 8'b11001000) ? {26'b10001111100011111101011110} :
                        (ma[22:15] == 8'b11001001) ? {26'b10001111001111111000001010} :
                        (ma[22:15] == 8'b11001010) ? {26'b10001110111011111000011101} :
                        (ma[22:15] == 8'b11001011) ? {26'b10001110100111111110010101} :
                        (ma[22:15] == 8'b11001100) ? {26'b10001110010100001001101110} :
                        (ma[22:15] == 8'b11001101) ? {26'b10001110000000011010101000} :
                        (ma[22:15] == 8'b11001110) ? {26'b10001101101100110000111111} :
                        (ma[22:15] == 8'b11001111) ? {26'b10001101011001001100110001} :
                        (ma[22:15] == 8'b11010000) ? {26'b10001101000101101101111100} :
                        (ma[22:15] == 8'b11010001) ? {26'b10001100110010010100011111} :
                        (ma[22:15] == 8'b11010010) ? {26'b10001100011111000000010101} :
                        (ma[22:15] == 8'b11010011) ? {26'b10001100001011110001011111} :
                        (ma[22:15] == 8'b11010100) ? {26'b10001011111000100111111000} :
                        (ma[22:15] == 8'b11010101) ? {26'b10001011100101100011100000} :
                        (ma[22:15] == 8'b11010110) ? {26'b10001011010010100100010100} :
                        (ma[22:15] == 8'b11010111) ? {26'b10001010111111101010010010} :
                        (ma[22:15] == 8'b11011000) ? {26'b10001010101100110101010111} :
                        (ma[22:15] == 8'b11011001) ? {26'b10001010011010000101100010} :
                        (ma[22:15] == 8'b11011010) ? {26'b10001010000111011010110001} :
                        (ma[22:15] == 8'b11011011) ? {26'b10001001110100110101000001} :
                        (ma[22:15] == 8'b11011100) ? {26'b10001001100010010100010001} :
                        (ma[22:15] == 8'b11011101) ? {26'b10001001001111111000011111} :
                        (ma[22:15] == 8'b11011110) ? {26'b10001000111101100001101000} :
                        (ma[22:15] == 8'b11011111) ? {26'b10001000101011001111101011} :
                        (ma[22:15] == 8'b11100000) ? {26'b10001000011001000010100110} :
                        (ma[22:15] == 8'b11100001) ? {26'b10001000000110111010010110} :
                        (ma[22:15] == 8'b11100010) ? {26'b10000111110100110110111010} :
                        (ma[22:15] == 8'b11100011) ? {26'b10000111100010111000010000} :
                        (ma[22:15] == 8'b11100100) ? {26'b10000111010000111110010110} :
                        (ma[22:15] == 8'b11100101) ? {26'b10000110111111001001001010} :
                        (ma[22:15] == 8'b11100110) ? {26'b10000110101101011000101010} :
                        (ma[22:15] == 8'b11100111) ? {26'b10000110011011101100110101} :
                        (ma[22:15] == 8'b11101000) ? {26'b10000110001010000101101000} :
                        (ma[22:15] == 8'b11101001) ? {26'b10000101111000100011000010} :
                        (ma[22:15] == 8'b11101010) ? {26'b10000101100111000101000001} :
                        (ma[22:15] == 8'b11101011) ? {26'b10000101010101101011100011} :
                        (ma[22:15] == 8'b11101100) ? {26'b10000101000100010110100111} :
                        (ma[22:15] == 8'b11101101) ? {26'b10000100110011000110001010} :
                        (ma[22:15] == 8'b11101110) ? {26'b10000100100001111010001011} :
                        (ma[22:15] == 8'b11101111) ? {26'b10000100010000110010101000} :
                        (ma[22:15] == 8'b11110000) ? {26'b10000011111111101111100000} :
                        (ma[22:15] == 8'b11110001) ? {26'b10000011101110110000110000} :
                        (ma[22:15] == 8'b11110010) ? {26'b10000011011101110110010111} :
                        (ma[22:15] == 8'b11110011) ? {26'b10000011001101000000010100} :
                        (ma[22:15] == 8'b11110100) ? {26'b10000010111100001110100100} :
                        (ma[22:15] == 8'b11110101) ? {26'b10000010101011100001000111} :
                        (ma[22:15] == 8'b11110110) ? {26'b10000010011010110111111010} :
                        (ma[22:15] == 8'b11110111) ? {26'b10000010001010010010111100} :
                        (ma[22:15] == 8'b11111000) ? {26'b10000001111001110010001011} :
                        (ma[22:15] == 8'b11111001) ? {26'b10000001101001010101100101} :
                        (ma[22:15] == 8'b11111010) ? {26'b10000001011000111101001010} :
                        (ma[22:15] == 8'b11111011) ? {26'b10000001001000101000110110} :
                        (ma[22:15] == 8'b11111100) ? {26'b10000000111000011000101010} :
                        (ma[22:15] == 8'b11111101) ? {26'b10000000101000001100100011} :
                        (ma[22:15] == 8'b11111110) ? {26'b10000000011000000100100000} : {26'b10000000001000000000100000};

   wire [25:0] x_out1;
   wire [25:0] x_out2;
   newton_inv u1(ma,x_out0,x_out1);
   newton_inv u2(ma,x_out1,x_out2);

   wire [22:0] my = (e == 8'd254) ? ((x_out2[3:3]) ? {1'b0,x_out2[25:4]} + 23'b1 : {1'b0,x_out2[25:4]}) :
                    (e == 8'd253) ? ((x_out2[2:2]) ? x_out2[25:3] + 23'b1 : x_out2[25:3]) :
                    (x_out2[1:1]) ? x_out2[24:2] + 23'b1 : x_out2[24:2];

   wire [7:0] ey = (e == 8'd254) ? 0 : 8'd253 - e;
   wire [7:0] ey2 = (e == 8'd253) ? 0 : ey + 8'b1;

   // nanかどうかの判定
   wire nzm = |x[22:0];
   assign y = (e == 8'd255 && nzm) ? {s,8'd255,1'b1,x[21:0]} : // 元がnanなら結果もnan
              (e == 8'd255 && ~nzm) ? {s,8'd0,23'b0} : // 元がinfなら結果は0
              (~|x) ? {s,8'd255,23'b0} : // 元が+-0なら結果は+-inf
              (~|x[22:0]) ? ((e == 8'd254) ? {s,8'b0,1'b1,22'b0} : (e == 8'd253) ? {s,8'b1,23'b0} : {s,ey2,23'b0}) : {s,ey,my};

   assign exception = (e == 8'd255 && nzm) ? 1'b1 : 1'b0;

endmodule

module fdiv
   (  input wire [31:0]  x1,
      input wire [31:0]  x2,
      output wire [31:0] y,
      output wire        ovf);
   // 定義
   wire s1 = x1[31:31];
   wire [7:0] e1 = x1[30:23];
   wire [22:0] m1 = x1[22:0];
   wire s2 = x2[31:31];
   wire [7:0] e2 = x2[30:23];
   wire [22:0] m2 = x2[22:0];
   // 非正規化数の処理
   // wire [23:0] m2a = (|e2) ? {1'b1,m2} :
   //                   (m2a[22:22]) ? {m2a[22:0],1'b0} :
   //                   (m2a[21:21]) ? {m2a[21:0],2'b0} :
   //                   (m2a[20:20]) ? {m2a[20:0],3'b0} :
   //                   (m2a[19:19]) ? {m2a[19:0],4'b0} :
   //                   (m2a[18:18]) ? {m2a[18:0],5'b0} :
   //                   (m2a[17:17]) ? {m2a[17:0],6'b0} :
   //                   (m2a[16:16]) ? {m2a[16:0],7'b0} :
   //                   (m2a[15:15]) ? {m2a[15:0],8'b0} :
   //                   (m2a[14:14]) ? {m2a[14:0],9'b0} :
   //                   (m2a[13:13]) ? {m2a[13:0],10'b0} :
   //                   (m2a[12:12]) ? {m2a[12:0],11'b0} :
   //                   (m2a[11:11]) ? {m2a[11:0],12'b0} :
   //                   (m2a[10:10]) ? {m2a[10:0],13'b0} :
   //                   (m2a[9:9]) ? {m2a[9:0],14'b0} :
   //                   (m2a[8:8]) ? {m2a[8:0],15'b0} :
   //                   (m2a[7:7]) ? {m2a[7:0],16'b0} :
   //                   (m2a[6:6]) ? {m2a[6:0],17'b0} :
   //                   (m2a[5:5]) ? {m2a[5:0],18'b0} :
   //                   (m2a[4:4]) ? {m2a[4:0],19'b0} :
   //                   (m2a[3:3]) ? {m2a[3:0],20'b0} :
   //                   (m2a[2:2]) ? {m2a[2:0],21'b0} :
   //                   (m2a[1:1]) ? {m2a[1:0],22'b0} : {m2a[0:0],23'b0};

   // wire [4:0] ee1 = (|e1) ? 5'd0 :
   //                 (m1a[22:22]) ? 5'd1 :
   //                 (m1a[21:21]) ? 5'd2 :
   //                 (m1a[20:20]) ? 5'd3 :
   //                 (m1a[19:19]) ? 5'd4 :
   //                 (m1a[18:18]) ? 5'd5 :
   //                 (m1a[17:17]) ? 5'd6 :
   //                 (m1a[16:16]) ? 5'd7 :
   //                 (m1a[15:15]) ? 5'd8 :
   //                 (m1a[14:14]) ? 5'd9 :
   //                 (m1a[13:13]) ? 5'd10 :
   //                 (m1a[12:12]) ? 5'd11 :
   //                 (m1a[11:11]) ? 5'd12 :
   //                 (m1a[10:10]) ? 5'd13 :
   //                 (m1a[9:9]) ? 5'd14 :
   //                 (m1a[8:8]) ? 5'd15 :
   //                 (m1a[7:7]) ? 5'd16 :
   //                 (m1a[6:6]) ? 5'd17 :
   //                 (m1a[5:5]) ? 5'd18 :
   //                 (m1a[4:4]) ? 5'd19 :
   //                 (m1a[3:3]) ? 5'd20 :
   //                 (m1a[2:2]) ? 5'd21 :
   //                 (m1a[1:1]) ? 5'd22 : 5'd23;
   // wire [4:0] ee2 = (|e2) ? 5'd0 :
   //                 (m2a[22:22]) ? 5'd1 :
   //                 (m2a[21:21]) ? 5'd2 :
   //                 (m2a[20:20]) ? 5'd3 :
   //                 (m2a[19:19]) ? 5'd4 :
   //                 (m2a[18:18]) ? 5'd5 :
   //                 (m2a[17:17]) ? 5'd6 :
   //                 (m2a[16:16]) ? 5'd7 :
   //                 (m2a[15:15]) ? 5'd8 :
   //                 (m2a[14:14]) ? 5'd9 :
   //                 (m2a[13:13]) ? 5'd10 :
   //                 (m2a[12:12]) ? 5'd11 :
   //                 (m2a[11:11]) ? 5'd12 :
   //                 (m2a[10:10]) ? 5'd13 :
   //                 (m2a[9:9]) ? 5'd14 :
   //                 (m2a[8:8]) ? 5'd15 :
   //                 (m2a[7:7]) ? 5'd16 :
   //                 (m2a[6:6]) ? 5'd17 :
   //                 (m2a[5:5]) ? 5'd18 :
   //                 (m2a[4:4]) ? 5'd19 :
   //                 (m2a[3:3]) ? 5'd20 :
   //                 (m2a[2:2]) ? 5'd21 :
   //                 (m2a[1:1]) ? 5'd22 : 5'd23;
                   
   // wire [5:0] edif = ee2 - ee1;

   // wire [45:0] mm = (e == 5'd0) ? {23'd0,m1} :
   //                   (e == 5'd1) ? {22'd0,m1,1'd0} :
   //                   (e == 5'd2) ? {21'd0,m1,2'd0} :
   //                   (e == 5'd3) ? {20'd0,m1,3'd0} :
   //                   (e == 5'd4) ? {19'd0,m1,4'd0} :
   //                   (e == 5'd5) ? {18'd0,m1,5'd0} :
   //                   (e == 5'd6) ? {17'd0,m1,6'd0} :
   //                   (e == 5'd7) ? {16'd0,m1,7'd0} :
   //                   (e == 5'd8) ? {15'd0,m1,8'd0} :
   //                   (e == 5'd9) ? {14'd0,m1,9'd0} :
   //                   (e == 5'd10) ? {13'd0,m1,10'd0} :
   //                   (e == 5'd11) ? {12'd0,m1,11'd0} :
   //                   (e == 5'd12) ? {11'd0,m1,12'd0} :
   //                   (e == 5'd13) ? {10'd0,m1,13'd0} :
   //                   (e == 5'd14) ? {9'd0,m1,14'd0} :
   //                   (e == 5'd15) ? {8'd0,m1,15'd0} :
   //                   (e == 5'd16) ? {7'd0,m1,16'd0} :
   //                   (e == 5'd17) ? {6'd0,m1,17'd0} :
   //                   (e == 5'd18) ? {5'd0,m1,18'd0} :
   //                   (e == 5'd19) ? {4'd0,m1,19'd0} :
   //                   (e == 5'd20) ? {3'd0,m1,20'd0} :
   //                   (e == 5'd21) ? {2'd0,m1,21'd0} :
   //                   (e == 5'd22) ? {1'd0,m1,22'd0} :
   //                   (e == 5'd23) ? {m1,23'd0} :

   // wire [22:0] m1a = (|e1) ? m1 :


   
   // wire [8:0] e1a = (|e1 && |e2) ? e1 :
   //                  (|e2) ? 8'b1 :
   //                  (|e1 && ~|e2) ?
   //                  ((m2a[22:22]) ? {1'b0,e1} + {9'd1} :
   //                   (m2a[21:21]) ? {1'b0,e1} + {9'd2} :
   //                   (m2a[20:20]) ? {1'b0,e1} + {9'd3} :
   //                   (m2a[19:19]) ? {1'b0,e1} + {9'd4} :
   //                   (m2a[18:18]) ? {1'b0,e1} + {9'd5} :
   //                   (m2a[17:17]) ? {1'b0,e1} + {9'd6} :
   //                   (m2a[16:16]) ? {1'b0,e1} + {9'd7} :
   //                   (m2a[15:15]) ? {1'b0,e1} + {9'd8} :
   //                   (m2a[14:14]) ? {1'b0,e1} + {9'd9} :
   //                   (m2a[13:13]) ? {1'b0,e1} + {9'd10} :
   //                   (m2a[12:12]) ? {1'b0,e1} + {9'd11} :
   //                   (m2a[11:11]) ? {1'b0,e1} + {9'd12} :
   //                   (m2a[10:10]) ? {1'b0,e1} + {9'd13} :
   //                   (m2a[9:9]) ? {1'b0,e1} + {9'd14} :
   //                   (m2a[8:8]) ? {1'b0,e1} + {9'd15} :
   //                   (m2a[7:7]) ? {1'b0,e1} + {9'd16} :
   //                   (m2a[6:6]) ? {1'b0,e1} + {9'd17} :
   //                   (m2a[5:5]) ? {1'b0,e1} + {9'd18} :
   //                   (m2a[4:4]) ? {1'b0,e1} + {9'd19} :
   //                   (m2a[3:3]) ? {1'b0,e1} + {9'd20} :
   //                   (m2a[2:2]) ? {1'b0,e1} + {9'd21} :
   //                   (m2a[1:1]) ? {1'b0,e1} + {9'd22} : {1'b0,e1} + {9'd23}) :
   //                  ((m2a[22:22]) ? {1'b0,e1} + {9'd2} :
   //                   (m2a[21:21]) ? {1'b0,e1} + {9'd3} :
   //                   (m2a[20:20]) ? {1'b0,e1} + {9'd4} :
   //                   (m2a[19:19]) ? {1'b0,e1} + {9'd5} :
   //                   (m2a[18:18]) ? {1'b0,e1} + {9'd6} :
   //                   (m2a[17:17]) ? {1'b0,e1} + {9'd7} :
   //                   (m2a[16:16]) ? {1'b0,e1} + {9'd8} :
   //                   (m2a[15:15]) ? {1'b0,e1} + {9'd9} :
   //                   (m2a[14:14]) ? {1'b0,e1} + {9'd10} :
   //                   (m2a[13:13]) ? {1'b0,e1} + {9'd11} :
   //                   (m2a[12:12]) ? {1'b0,e1} + {9'd12} :
   //                   (m2a[11:11]) ? {1'b0,e1} + {9'd13} :
   //                   (m2a[10:10]) ? {1'b0,e1} + {9'd14} :
   //                   (m2a[9:9]) ? {1'b0,e1} + {9'd15} :
   //                   (m2a[8:8]) ? {1'b0,e1} + {9'd16} :
   //                   (m2a[7:7]) ? {1'b0,e1} + {9'd17} :
   //                   (m2a[6:6]) ? {1'b0,e1} + {9'd18} :
   //                   (m2a[5:5]) ? {1'b0,e1} + {9'd19} :
   //                   (m2a[4:4]) ? {1'b0,e1} + {9'd20} :
   //                   (m2a[3:3]) ? {1'b0,e1} + {9'd21} :
   //                   (m2a[2:2]) ? {1'b0,e1} + {9'd22} :
   //                   (m2a[1:1]) ? {1'b0,e1} + {9'd23} : {1'b0,e1} + {9'd24});

   // wire [7:0] e2a = (|e2) ? e2 : 8'b1;

   wire [31:0] x2i;
   wire exception;
   finv u1(x2,x2i,exception);

   // wire ex;
   wire [31:0] my;
   fmul u2(x2i,x1,my,ovf);

   assign y = my;
   // assign ovf = (e1a[8:8] || ex) ? 1'b1 : 1'b0;

endmodule                                                                         
`default_nettype wire